library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom_bcd is
    port (
		  clock : in std_logic;
        dataout : out std_logic_vector (11 downto 0);
        address : in std_logic_vector (7 downto 0)
    );
end entity;

architecture arch of rom_bcd is

    subtype word is std_logic_vector (11 downto 0);
    type word_array is array (255 downto 0) of word;

    constant memory : word_array := (
			x"255",
			x"254",
			x"253",
			x"252",
			x"251",
			x"250",
			x"249",
			x"248",
			x"247",
			x"246",
			x"245",
			x"244",
			x"243",
			x"242",
			x"241",
			x"240",
			x"239",
			x"238",
			x"237",
			x"236",
			x"235",
			x"234",
			x"233",
			x"232",
			x"231",
			x"230",
			x"229",
			x"228",
			x"227",
			x"226",
			x"225",
			x"224",
			x"223",
			x"222",
			x"221",
			x"220",
			x"219",
			x"218",
			x"217",
			x"216",
			x"215",
			x"214",
			x"213",
			x"212",
			x"211",
			x"210",
			x"209",
			x"208",
			x"207",
			x"206",
			x"205",
			x"204",
			x"203",
			x"202",
			x"201",
			x"200",
			x"199",
			x"198",
			x"197",
			x"196",
			x"195",
			x"194",
			x"193",
			x"192",
			x"191",
			x"190",
			x"189",
			x"188",
			x"187",
			x"186",
			x"185",
			x"184",
			x"183",
			x"182",
			x"181",
			x"180",
			x"179",
			x"178",
			x"177",
			x"176",
			x"175",
			x"174",
			x"173",
			x"172",
			x"171",
			x"170",
			x"169",
			x"168",
			x"167",
			x"166",
			x"165",
			x"164",
			x"163",
			x"162",
			x"161",
			x"160",
			x"159",
			x"158",
			x"157",
			x"156",
			x"155",
			x"154",
			x"153",
			x"152",
			x"151",
			x"150",
			x"149",
			x"148",
			x"147",
			x"146",
			x"145",
			x"144",
			x"143",
			x"142",
			x"141",
			x"140",
			x"139",
			x"138",
			x"137",
			x"136",
			x"135",
			x"134",
			x"133",
			x"132",
			x"131",
			x"130",
			x"129",
			x"128",
			x"127",
			x"126",
			x"125",
			x"124",
			x"123",
			x"122",
			x"121",
			x"120",
			x"119",
			x"118",
			x"117",
			x"116",
			x"115",
			x"114",
			x"113",
			x"112",
			x"111",
			x"110",
			x"109",
			x"108",
			x"107",
			x"106",
			x"105",
			x"104",
			x"103",
			x"102",
			x"101",
			x"100",
			x"099",
			x"098",
			x"097",
			x"096",
			x"095",
			x"094",
			x"093",
			x"092",
			x"091",
			x"090",
			x"089",
			x"088",
			x"087",
			x"086",
			x"085",
			x"084",
			x"083",
			x"082",
			x"081",
			x"080",
			x"079",
			x"078",
			x"077",
			x"076",
			x"075",
			x"074",
			x"073",
			x"072",
			x"071",
			x"070",
			x"069",
			x"068",
			x"067",
			x"066",
			x"065",
			x"064",
			x"063",
			x"062",
			x"061",
			x"060",
			x"059",
			x"058",
			x"057",
			x"056",
			x"055",
			x"054",
			x"053",
			x"052",
			x"051",
			x"050",
			x"049",
			x"048",
			x"047",
			x"046",
			x"045",
			x"044",
			x"043",
			x"042",
			x"041",
			x"040",
			x"039",
			x"038",
			x"037",
			x"036",
			x"035",
			x"034",
			x"033",
			x"032",
			x"031",
			x"030",
			x"029",
			x"028",
			x"027",
			x"026",
			x"025",
			x"024",
			x"023",
			x"022",
			x"021",
			x"020",
			x"019",
			x"018",
			x"017",
			x"016",
			x"015",
			x"014",
			x"013",
			x"012",
			x"011",
			x"010",
			x"009",
			x"008",
			x"007",
			x"006",
			x"005",
			x"004",
			x"003",
			x"002",
			x"001",
			x"000"
   );

begin
		sync: process (clock)
			begin
			  if rising_edge(clock) then
				 dataout <= memory(to_integer(unsigned(address)));
			  end if;
			end process sync;
      
end architecture;
